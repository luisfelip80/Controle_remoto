module ula(clock,a,b,r,op,sb,sa,enable,sinA, sinB);
	input [7:0]a;
	input [7:0]b;
	input op;
	input clock;
	output reg [8:0]r;
	output sa, sb;
	input sinA;
	input sinB;
	reg saa;
	reg sbb;
	reg sinal;
	input enable;
	reg [6:0]aa;
	reg [6:0]bb;
	reg [7:0]rr;
	always @(posedge clock) begin
		saa = sinA;
		sbb = sinB;
		aa = a[6:0];
		bb = b[6:0];
		case(op)
			0: begin
				if(saa == 0 && sbb == 0)begin
					rr = aa + bb;
					sinal = 0;
				end
				if(saa == 1 && sbb == 0)begin
					if(aa > bb)begin
						rr = aa - bb;
						sinal = saa;
					end
					else begin
						rr = bb - aa;
						sinal = sbb;
					end
				end
				if(saa == 0 && sbb == 1)begin
					if(aa > bb)begin
						rr = aa - bb;
						sinal = saa;
					end
					else begin
						rr = bb - aa;
						sinal = sbb;
					end
				end
				if(saa == 1 && sbb == 1)begin
					rr = aa + bb;
					sinal = 1;
				end
			end	
			1: begin
			sbb = ~sbb;
			if(saa == 0 && sbb == 0)begin
					rr = aa + bb;
					sinal = 0;
				end
				if(saa == 1 && sbb == 0)begin
					if(aa > bb)begin
						rr = aa - bb;
						sinal = saa;
					end
					else begin
						rr = bb - aa;
						sinal = sbb;
					end
				end
				if(saa == 0 && sbb == 1)begin
					if(aa > bb)begin
						rr = aa - bb;
						sinal = saa;
					end
					else begin
						rr = bb - aa;
						sinal = sbb;
					end
				end
				if(saa == 1 && sbb == 1)begin
					rr = aa + bb;
					sinal = 1;
				end
			end	
		endcase

	end
	always @(posedge clock) begin
		if (rr==0) begin
			r[8] <= 1;
			r[7:0] = rr;
		end
		else begin
			r[8] <= ~sinal;
			r[7:0] = rr;
		end
	end
	assign sa = saa;
	assign sb = sbb;


endmodule