module up_counter(out,enable,clk,reset);
  output reg [16:0] out;
  input enable;
  input clk;
  input reset;  
  //-------------Code Starts Here-------
  always @(posedge clk)begin
  	if (reset) begin
  		out <= 0 ;
  	end 
  	else if (enable) begin
  		out <= out + 1;
  	end
	
  end
endmodule
