module Remoto (comando,comparador,clk,entrada,led);
	output reg [7:0] comando;
	output reg [7:0]comparador;
	input clk;
	input entrada;
	output reg led;
	reg [7:0]cont;
	reg [7:0]etapa;
	reg enable,reset,b,enableO;
	reg [7:0]bitSgnal;
	wire [16:0]tempoWire;
	wire [7:0]copia1;
	reg [7:0]copia2;
	reg [16:0]tempo;
	initial begin
		led = 0;
		etapa = 0;
		enable = 0;
		comando =0;
		cont = 0;
		reset = 0;
		b = 0;
		bitSgnal = 0;
	end
	up_counter G2(.out(tempoWire),.enable(enable),.clk(clk),.reset(reset));
	orgBits G1(.ordem(bitSgnal),.b(b),.out(copia1),.in(copia2),.clk(clk),.enable(enableO));

	always@(posedge clk)begin
		
		if(entrada==0 && etapa==0)begin
			etapa <= 1;
			enable<= 1;
			reset <=0;
			tempo <= 0;
		end
		if(entrada==1 && etapa == 1)begin
			tempo <= tempoWire;
			enable<= 0;
			reset <=1;
			if (tempo > 23000)begin
				tempo <= 0;
				etapa <=2;
				enable<= 0;
				reset <=1;
				if(led)begin
					led<=0;
				end
				else begin
					led<=1;
				end
			end
			tempo <= 0;
		end
		if(entrada==0 && etapa == 2 )begin
			etapa <= 3;
			if(cont == 16)begin
				cont <= 0;
				etapa <= 4;
			end
		end
		if(entrada == 1 && etapa == 3)begin
			etapa <= 2;
			cont <= cont + 1;
		end
		if(entrada ==1 && etapa == 4)begin
			enable<= 1;
			etapa <= 5;
			reset <=0;
			cont <= cont + 1;
		end 
		else if(entrada == 0 && etapa == 5)begin
			enable <=0;
			reset <=1;
			if(cont == 8) begin
				cont <= 0;
				etapa <=6;
				bitSgnal <= 0;
				comando = copia2;
				reset <= 0;
			end
			else begin 
				etapa <=4;
			end
			tempo <= tempoWire;
			if(tempo > 23000)begin // bit = 1 
				tempo <= 0;
				b<= 1;
				copia2 <= copia1;
				enableO <= 0;
				bitSgnal <= bitSgnal + 1;
				enableO<=1;
				if(bitSgnal==8)begin
					bitSgnal <= 0;
				end
			end
			else if (tempo <= 23000)begin// bit = 0
				b<= 0;
				tempo <= 0;
				enableO <= 1;
				copia2 <= copia1;
				enableO <= 0;
				bitSgnal <= bitSgnal + 1;
				if(bitSgnal==8)begin
					bitSgnal <= 0;
				end
			end
		end
		
		if(entrada == 1 && etapa == 6)begin
			enable<= 1;
			etapa <= 7;
			reset <=0;
			cont <= cont + 1;
		end 
		else if(entrada == 0 && etapa == 7)begin
			enable <=0;
			reset <=1;
			if(cont == 8) begin
				cont <= 0;
				etapa <=8;
				bitSgnal <= 0;
				comparador <= copia2;
				reset <= 0;
			end
			else begin
				etapa <=6;
			end
			tempo<=tempoWire;
			if(tempo > 23000)begin // bit = 1 
				tempo <= 0;
				b <= 1;
				//orgBits(.ordem(bitSgnal),.b(b),.out(copia),.clk(clk));
				enableO <= 1;
				copia2 <= copia1;
				enableO <= 0;
				bitSgnal <= bitSgnal + 1;
				if(bitSgnal==8)begin
					bitSgnal <= 0;
				end
			end
			else if (tempo <= 23000)begin// bit = 0
				tempo <= 0;
				b<= 0;
				enableO <= 1;
				copia2 <= copia1;
				enableO <= 0;
				//orgBits(.ordem(bitSgnal),.b(b),.out(copia),.clk(clk));
				bitSgnal <= bitSgnal + 1;
				if(bitSgnal==8)begin
					bitSgnal <= 0;
				end
			end
		end
		if(etapa==8) begin
			cont <= 0;
			etapa <=0;
			bitSgnal <= 0;
			reset <= 0;
			tempo <= 0;
		end
	end
endmodule
